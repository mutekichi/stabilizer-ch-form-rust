0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,-1.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
0.000000000000000000e+00,0.000000000000000000e+00
