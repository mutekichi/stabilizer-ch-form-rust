2.077481888934145469e-17,-6.980756726287458820e-18
-1.125016984820677569e-17,-5.501801922474044400e-18
1.249999999999991396e-01,1.249999999999991118e-01
-7.653810781896326339e-18,-1.113051595930492550e-17
2.832321140486134431e-18,-8.171282704461957450e-18
-3.469446951953613418e-18,5.501801922474044400e-18
1.249999999999991812e-01,1.249999999999991535e-01
-1.256034971528312296e-17,9.686165752416756550e-18
9.771215044393362809e-18,1.679383459306105207e-17
2.627617959607677601e-18,-1.437091981433183015e-18
1.249999999999991257e-01,-1.249999999999991396e-01
1.400469992217129192e-17,1.891123885555808854e-17
-1.104546666732832232e-17,-9.771215044393362809e-18
1.818906375211400407e-17,1.328252481872720744e-17
1.249999999999991396e-01,-1.249999999999991535e-01
2.094359382607851721e-17,-2.747271848509529328e-18
-9.854940689153823693e-18,-3.761051630478273720e-17
-3.469446951953613804e-18,8.418289923459350475e-19
-1.249999999999991396e-01,-1.249999999999991535e-01
-1.256034971528312296e-17,1.112325773384993899e-17
-1.958429291116695606e-17,4.186282238023044213e-20
5.501801922474043630e-18,2.250033969641355138e-17
1.249999999999991673e-01,1.249999999999991396e-01
1.746688864866991959e-17,2.728722474089849627e-17
-1.679383459306105207e-17,-1.671010894830059119e-17
3.900574546383568612e-17,1.100360384494808880e-17
-1.249999999999991673e-01,1.249999999999991535e-01
1.269121143568363161e-19,-7.149168779890988277e-19
-4.733986852679586957e-17,1.671010894830059119e-17
-2.106324771498036894e-17,3.469446951953613418e-18
1.249999999999991535e-01,-1.249999999999991535e-01
-1.113051595930492550e-17,1.399744169671630540e-17
3.589100840855465146e-18,7.653810781896326339e-18
-1.249999999999991535e-01,1.249999999999991396e-01
-8.375985885340410814e-18,-1.437091981433183207e-18
6.980756726287458820e-18,-1.679383459306105207e-17
-1.400469992217129192e-17,-3.001096077223203116e-18
-1.249999999999991535e-01,1.249999999999991535e-01
-5.952629890872474856e-19,3.469446951953613418e-18
-1.671010894830059119e-17,1.958429291116695606e-17
-2.296869057114396553e-17,1.746688864866991959e-17
1.249999999999991396e-01,1.249999999999991396e-01
-1.531487978924763611e-17,2.165851070406761825e-17
-6.980756726287458820e-18,2.832321140486134431e-18
-2.356395356023121176e-17,6.216718800463143902e-18
1.249999999999991535e-01,1.249999999999991396e-01
-4.906538933386798166e-18,-6.343630914819979833e-18
2.652318681507418444e-17,9.771215044393362809e-18
3.589100840855465146e-18,-2.159267084877267298e-18
1.249999999999991535e-01,-1.249999999999991257e-01
-4.311275944299548851e-18,-8.583538376948312719e-35
-1.671010894830059119e-17,2.652318681507418444e-17
-9.686165752416756550e-18,1.256760794073810794e-17
-1.249999999999991535e-01,1.249999999999991396e-01
2.716031262654166111e-17,2.141194470080892829e-17
-4.186282238023044213e-20,2.779743843800914395e-17
2.754530073964515072e-18,-6.223977025918128876e-18
-1.249999999999991673e-01,-1.249999999999991673e-01
1.209199884055271189e-17,-1.962615573354718650e-17
2.939737077794054931e-17,-4.186282238023044213e-20
-6.223977025918128105e-18,-1.399744169671630540e-17
1.249999999999991257e-01,1.249999999999991535e-01
-1.387778780781445367e-17,2.309560268550080069e-17
9.854940689153823693e-18,2.660691245983464532e-17
5.621455811375896127e-18,-4.184363829942713691e-18
-1.249999999999990979e-01,-1.249999999999991396e-01
-1.437091981433183207e-18,6.938893903907226067e-18
-3.058789675611504794e-17,2.660691245983464532e-17
5.621455811375895357e-18,2.931957971141892494e-17
-1.249999999999991673e-01,-1.249999999999991673e-01
1.531487978924763919e-17,-2.369086567458805001e-17
2.204907051227641421e-17,3.067162240087550883e-17
-1.891123885555808854e-17,1.375087569345761697e-17
-1.249999999999991673e-01,1.249999999999991396e-01
-1.447305079690169991e-17,1.065490685911952945e-17
1.104546666732832232e-17,2.832321140486134431e-18
-2.991484270050617426e-17,-7.661069007351311313e-18
-1.249999999999991257e-01,1.249999999999991396e-01
2.022141872263443274e-17,-8.375985885340410814e-18
9.854940689153823693e-18,-3.067162240087550883e-17
5.621455811375895357e-18,1.459996291125853815e-17
1.249999999999991535e-01,1.249999999999991257e-01
1.184543283729402346e-17,2.410663727404873470e-34
-2.832321140486134431e-18,6.980756726287458820e-18
-1.028142874150400432e-17,-9.693423977871741524e-18
-1.249999999999991396e-01,-1.249999999999991535e-01
-5.501801922474044400e-18,1.591014277833488543e-17
-1.679383459306105207e-17,1.264539900725972768e-17
-2.381777778894488517e-17,5.374889808117206928e-18
1.249999999999991535e-01,-1.249999999999991396e-01
8.375985885340409274e-18,-6.938893903907226067e-18
-1.958429291116695606e-17,1.264539900725972768e-17
2.788248772998574559e-17,3.625847361532615949e-17
-1.249999999999991396e-01,1.249999999999991257e-01
-9.566511863514904823e-18,2.874183962866365644e-18
1.671010894830059119e-17,-2.832321140486134431e-18
-4.186282238023044213e-20,4.186282238023044213e-20
-8.971248874427658589e-18,-1.100360384494808880e-17
1.249999999999991673e-01,-1.249999999999991396e-01
2.991484270050617426e-17,2.644539574855256315e-17
-9.854940689153823693e-18,-9.771215044393362809e-18
7.534156892994474611e-18,-4.064709941040860423e-18
1.249999999999991535e-01,-1.249999999999991535e-01
-7.407244778637637910e-18,-2.787522950453076216e-17
-2.832321140486134431e-18,1.232388800554729073e-18
-2.874183962866364874e-18,2.943923360032077975e-17
-1.249999999999991673e-01,-1.249999999999991535e-01
-2.034833083699127098e-17,3.422611864480572465e-17
-3.058789675611504794e-17,-4.040097462288864119e-17
-4.906538933386796626e-18,1.184543283729402192e-17
-1.249999999999991396e-01,-1.249999999999991118e-01
3.074941346739712703e-17,5.628714036830881101e-18
1.671010894830059119e-17,-3.058789675611504794e-17
-1.962615573354718650e-17,-2.369086567458804693e-17
-1.249999999999991118e-01,1.249999999999991535e-01
7.065806018264063538e-18,3.278902666337254530e-17
1.232388800554729073e-18,-4.186282238023044213e-20
8.375985885340410814e-18,6.343630914819980603e-18
1.249999999999991535e-01,-1.249999999999991673e-01
-1.256760794073810948e-17,8.249073770983572572e-18
-3.633626468184777769e-17,-2.245847687403332093e-17
2.572322064510847868e-17,-1.675197177068082163e-17
1.249999999999991535e-01,1.249999999999991535e-01
1.806215163775716582e-17,7.065806018264065079e-18
-4.186282238023044213e-20,-6.980756726287458820e-18
-1.387778780781445367e-17,2.225377369315486449e-17
-1.249999999999991257e-01,-1.249999999999991118e-01
-9.090902763329508776e-18,-5.628714036830881872e-18
