1.864746193260806779e-17,-2.110010742601988100e-17
5.095193435455063994e-17,8.425799482132585271e-19
8.724994857809758860e-18,-1.573548229877980165e-17
-4.987079758440086470e-17,1.230276807527998464e-17
-2.439582985834080062e-17,1.434901683940504261e-17
-2.756764531575078399e-17,-1.200557554996287897e-17
-1.088083008963831695e-18,4.308510015434846504e-17
-2.661642711538013981e-17,-2.577397414975260464e-17
1.022041055598272537e-17,6.455775245048623534e-19
-2.329841962948503791e-19,1.633343449274248486e-18
-6.640950422722808857e-18,1.379092554799810177e-17
2.906969658207353350e-17,-1.371808406437210791e-17
4.593105756077906619e-17,-2.277606821603037579e-17
-1.224382038525861546e-17,-4.078915721286266098e-18
-2.009844770764587029e-17,-3.381621978537719874e-17
1.524578214531111551e-18,-3.362753852963175229e-17
-3.662544446335400271e-17,-1.025651931115494362e-17
2.088965017793338617e-17,-3.935306752051532956e-17
-1.366701857308717784e-17,1.235320959328333115e-17
-6.902473162094221433e-18,-2.754543035418322124e-17
-1.392810234323207451e-17,-9.676213058180421532e-18
-1.536519432466523846e-17,-4.431961708643159638e-17
-3.944130470948057888e-17,-2.596947466172635992e-17
-4.407198814066478691e-17,-5.137747792572477836e-20
-4.303359569383700674e-17,4.419633408480225293e-17
-1.754348622760914008e-17,-7.854315335746467668e-18
-2.148447419779411496e-17,1.752189523932312699e-17
3.621842376078564542e-17,1.790670098032389688e-17
-7.235774442583537645e-18,-3.335212199665572120e-17
-6.481119696694733574e-18,2.472062496681207875e-17
-5.153330355003328153e-17,-1.056742062602159707e-17
-5.684642421676189026e-17,4.529799890072990944e-17
8.838834764831762780e-02,-8.838834764831762780e-02
-8.838834764831760005e-02,8.838834764831758617e-02
-8.838834764831762780e-02,8.838834764831762780e-02
-8.838834764831762780e-02,8.838834764831760005e-02
8.838834764831762780e-02,8.838834764831760005e-02
8.838834764831758617e-02,8.838834764831762780e-02
8.838834764831762780e-02,8.838834764831760005e-02
-8.838834764831765556e-02,-8.838834764831760005e-02
8.838834764831762780e-02,-8.838834764831765556e-02
-8.838834764831762780e-02,8.838834764831761392e-02
-8.838834764831762780e-02,8.838834764831765556e-02
-8.838834764831757229e-02,8.838834764831762780e-02
-8.838834764831757229e-02,-8.838834764831762780e-02
-8.838834764831765556e-02,-8.838834764831762780e-02
-8.838834764831753066e-02,-8.838834764831761392e-02
8.838834764831762780e-02,8.838834764831762780e-02
8.838834764831762780e-02,8.838834764831764168e-02
-8.838834764831765556e-02,-8.838834764831761392e-02
-8.838834764831764168e-02,-8.838834764831766944e-02
-8.838834764831764168e-02,-8.838834764831757229e-02
8.838834764831765556e-02,-8.838834764831760005e-02
8.838834764831765556e-02,-8.838834764831761392e-02
8.838834764831762780e-02,-8.838834764831760005e-02
-8.838834764831764168e-02,8.838834764831762780e-02
-8.838834764831765556e-02,-8.838834764831761392e-02
8.838834764831765556e-02,8.838834764831760005e-02
8.838834764831764168e-02,8.838834764831764168e-02
8.838834764831766944e-02,8.838834764831764168e-02
8.838834764831757229e-02,-8.838834764831768331e-02
8.838834764831762780e-02,-8.838834764831764168e-02
8.838834764831760005e-02,-8.838834764831762780e-02
-8.838834764831764168e-02,8.838834764831757229e-02
2.700147456592872360e-18,-1.447273881026089734e-17
1.636685404303924918e-17,-6.205703163718680141e-18
-1.748305282940634600e-18,-7.043402104711703284e-19
2.215301763973388944e-17,1.709991780064204555e-17
-3.629126524441164698e-17,3.614193959283225022e-18
-6.641574396004393190e-18,-2.170926420871175346e-17
-4.884011985178428227e-18,7.668347616762208905e-17
3.062114262744475903e-18,5.009577259937357240e-17
1.463213056706244824e-17,-3.979682095153745938e-17
2.715104192705615381e-18,-2.619488864592557890e-17
-2.388774111571069346e-17,6.538224082813036943e-17
-1.432122925219578709e-17,-4.325481724544973786e-18
8.165216650613113412e-18,2.896756559950365180e-17
1.974912674853571814e-17,-2.724717488635799453e-17
-3.868558702108367149e-17,8.361780105095000517e-18
1.389136961477826500e-17,-3.716964196115629884e-17
-3.282181829245803895e-17,-2.474283992837966307e-17
-2.992585833725061953e-17,-3.718415972804251787e-17
7.730408360835546824e-18,-3.528835757947445989e-17
-9.914457893476151859e-18,2.748047106929364801e-17
-1.363090981791496422e-17,-6.256144681722035889e-18
-2.374161917923216980e-17,-3.977223707942915708e-18
2.965044180427456379e-17,7.470845337931593376e-19
-1.487975951282924230e-17,-8.774373433304984325e-18
1.142420635448024817e-17,5.923028405287815068e-18
1.272368257145295120e-17,6.379965088350026231e-17
3.641498721526750787e-17,4.000062642792101311e-18
4.979507399598513068e-18,6.540506355942630986e-18
4.355592456449043194e-19,-2.293652291534003695e-17
2.780632912027305180e-17,-5.025622729868323664e-17
-2.304528815008316445e-17,-8.774373433305005895e-18
1.487975951282925463e-17,-2.380056686925356363e-17
8.838834764831765556e-02,-8.838834764831758617e-02
-8.838834764831758617e-02,8.838834764831762780e-02
-8.838834764831762780e-02,8.838834764831760005e-02
-8.838834764831761392e-02,8.838834764831761392e-02
8.838834764831761392e-02,8.838834764831761392e-02
8.838834764831760005e-02,8.838834764831762780e-02
8.838834764831761392e-02,8.838834764831760005e-02
-8.838834764831762780e-02,-8.838834764831764168e-02
-8.838834764831768331e-02,8.838834764831762780e-02
8.838834764831765556e-02,-8.838834764831760005e-02
8.838834764831764168e-02,-8.838834764831764168e-02
8.838834764831766944e-02,-8.838834764831766944e-02
8.838834764831761392e-02,8.838834764831761392e-02
8.838834764831760005e-02,8.838834764831760005e-02
8.838834764831761392e-02,8.838834764831760005e-02
-8.838834764831762780e-02,-8.838834764831764168e-02
-8.838834764831761392e-02,-8.838834764831762780e-02
8.838834764831761392e-02,8.838834764831762780e-02
8.838834764831765556e-02,8.838834764831761392e-02
8.838834764831761392e-02,8.838834764831764168e-02
-8.838834764831760005e-02,8.838834764831762780e-02
-8.838834764831758617e-02,8.838834764831764168e-02
-8.838834764831758617e-02,8.838834764831762780e-02
8.838834764831764168e-02,-8.838834764831761392e-02
-8.838834764831761392e-02,-8.838834764831765556e-02
8.838834764831761392e-02,8.838834764831762780e-02
8.838834764831762780e-02,8.838834764831766944e-02
8.838834764831758617e-02,8.838834764831761392e-02
8.838834764831764168e-02,-8.838834764831758617e-02
8.838834764831762780e-02,-8.838834764831762780e-02
8.838834764831761392e-02,-8.838834764831758617e-02
-8.838834764831762780e-02,8.838834764831762780e-02
